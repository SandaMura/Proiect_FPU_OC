library verilog;
use verilog.vl_types.all;
entity test_log is
end test_log;
