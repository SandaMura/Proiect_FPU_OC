library verilog;
use verilog.vl_types.all;
entity testBench_adunare is
end testBench_adunare;
