library verilog;
use verilog.vl_types.all;
entity testBench_impartire is
end testBench_impartire;
