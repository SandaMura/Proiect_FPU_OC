library verilog;
use verilog.vl_types.all;
entity testBench_inmutire is
end testBench_inmutire;
